library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;  

entity SYED_Instruction is
port (
 SYED_Read_Address: in std_logic_vector(31 downto 0);
 SYED_Instruction: out  std_logic_vector(31 downto 0)
);
end SYED_Instruction;

architecture arch of SYED_Instruction is
signal SYED_ROM_Address: std_logic_vector(4 downto 0);
 type SYED_ROM_Type is array (0 to 31 ) of std_logic_vector(31 downto 0);
 constant SYED_ROM_Data: SYED_ROM_Type:=(
   "10001101010010000000000000000000",
	--100011 lw | 01010 register 10, 01000 dest. register , 0000 0000 offset, 0000
   "10001101011010010000000000000000", 
	--100011 lw | 01011 register 10, 01001 dest. register , 0000 0000 offset, 0000
   "10001101100010100000000000000000", 
	--100011 lw | 01100 register 10, 01010 dest. register , 0000 0000 offset, 0000
   "10001101101010110000000000000000", 
	--100011 lw | 01101 register 10, 01011 dest. register , 0000 0000 offset, 0000
   "10001111100011000000000000000000", 
	--100011 lw | 11100 register 10, 01100 dest. register , 0000 0000 offset, 0000
   "00000001000010011010100000000000", 
	--000000 add (R-type) | rs 01000 | rt 01001 | rd 10101
   "00000001010101011010100000000000", 
	--000000 add (R-type) | rs 01010 | rt 10101 | rd 10101
   "00000001011101011010100000000000", 
	--000000 add (R-type) | rs 01011 | rt 10101 | rd 10101
   "00000001100101011010100000000000",
	--000000 add (R-type) | rs 01100 | rt 10101 | rd 10101
   "10101101000100000000000000000000",
	--101011 sw | 01000 register 8, $t0 | 10000 register 16, $s0. $t0 = $s0
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
	"00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000",
   "00000000000000000000000000000000"
  );
begin

 SYED_ROM_Address <= SYED_Read_Address(5 downto 1);
  SYED_Instruction <= SYED_ROM_Data((to_integer(unsigned(SYED_ROM_Address)))/2) when SYED_Read_Address < x"00000020" else x"00000000";

end arch;